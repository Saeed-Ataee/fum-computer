//memory unit
module IMemBank(input memread, input [7:0] address, output reg [31:0] readdata);
 
  reg [31:0] mem_array [63:0];
  
  integer i;
  initial begin
      for (i=0; i<64; i=i+1)   
     mem_array[i]=i*10;
  end
 
  always@(memread, address, mem_array[address])begin
    if(memread)begin
      readdata=mem_array[address];
    end
  end

endmodule

module testbench;
  reg memread;              /* rw=RegWrite */
  reg [7:0] adr;  /* adr=address */
  wire [31:0] rd; /* rd=readdata */
  
  memBank u0(memread, adr, rd);
  
  initial begin
    memread=1'b0;
    adr=16'd0;
    
    #5
    memread=1'b1;
    adr=16'd0;
  end
  
  initial repeat(127)#4 adr=adr+1;
  
endmodule;
